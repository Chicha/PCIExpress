//======================================================
// Module name: key_test.v
// ����: ��⿪�����ϵ��ĸ�����KEY1~KEY4, ����⵽��������ʱ,��Ӧ��LED�Ʒ�ת
//======================================================
`timescale 1ns / 1ps
module key_test  (
							clk,              // ������������ʱ��: 100Mhz
							key_in,           // ���밴���ź�(KEY1~KEY4)
							led_out       // ���LED��,���ڿ��ƿ��������ĸ�LED(LED1~LED4)
						);

//========================================================
// PORT declarations
//========================================================						
input        clk; 
input  [1:0] key_in;
output [1:0] led_out;

wire rst_n=1'b1;

//�Ĵ�������
reg [19:0] count;
reg [1:0] key_scan; //����ɨ��ֵKEY

//==============================================
// ��������ֵ��20msɨ��һ��,����Ƶ��С�ڰ���ë��Ƶ�ʣ��൱���˳����˸�Ƶë���źš�
//==============================================
always @(posedge clk or negedge rst_n)     //���ʱ�ӵ������غ͸�λ���½���
begin
   if(!rst_n)                //��λ�źŵ���Ч
      count <= 20'd0;        //��������0
   else
      begin
         if(count ==20'd999_999)   //20msɨ��һ�ΰ���,20ms����(50M/50-1=999_999)
            begin
               count <= 20'b0;     //�������Ƶ�20ms������������
               key_scan <= key_in; //�������������ƽ
            end
         else
            count <= count + 20'b1; //��������1
     end
end
//====================================================
// �����ź�����һ��ʱ�ӽ���
//====================================================
reg [1:0] key_scan_r;
always @(posedge clk)
    key_scan_r <= key_scan;       
    
wire [1:0] flag_key = key_scan_r[1:0] & (~key_scan[1:0]);  //����⵽�������½��ر仯ʱ������ð��������£�������Ч 

//=====================================================
// LED�ƿ���,��������ʱ,��ص�LED�����ת
//=====================================================
reg [1:0] temp_led;
always @ (posedge clk or negedge rst_n)      //���ʱ�ӵ������غ͸�λ���½���
begin
    if (!rst_n)                 //��λ�źŵ���Ч
         temp_led <= 2'b11;   //LED�ƿ����ź����Ϊ��, LED��ȫ��
    else
         begin            
             if ( flag_key[0] ) temp_led[0] <= ~temp_led[0];   //����KEY1ֵ�仯ʱ��LED1��������ת
             if ( flag_key[1] ) temp_led[1] <= ~temp_led[1];   //����KEY2ֵ�仯ʱ��LED2��������ת
            
         end
end
 
 assign led_out[0] = temp_led[0];
 assign led_out[1] = temp_led[1];
 
            
endmodule
